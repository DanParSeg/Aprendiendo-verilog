//testbench for bf_cpu

module bf_cpu_tb();
    



endmodule